`define VERSION 007