module accelerator (arst_i,
    clk_i,
    done,
    start,
    data_in,
    data_out);
 input arst_i;
 input clk_i;
 output done;
 input start;
 input [31:0] data_in;
 output [31:0] data_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire clknet_0_clk_i;
 wire state;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_1_1__leaf_clk_i;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;

 sky130_fd_sc_hd__inv_2 _145_ (.A(net18),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _146_ (.A(net20),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _147_ (.A(net21),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _148_ (.A(net22),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _149_ (.A(net23),
    .Y(_118_));
 sky130_fd_sc_hd__inv_2 _150_ (.A(net25),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _151_ (.A(net48),
    .Y(_000_));
 sky130_fd_sc_hd__and2b_1 _152_ (.A_N(state),
    .B(net34),
    .X(_120_));
 sky130_fd_sc_hd__nor2_1 _153_ (.A(net73),
    .B(net47),
    .Y(_121_));
 sky130_fd_sc_hd__nand2_1 _154_ (.A(net8),
    .B(net31),
    .Y(_122_));
 sky130_fd_sc_hd__or2_1 _155_ (.A(net8),
    .B(net31),
    .X(_123_));
 sky130_fd_sc_hd__nand2_1 _156_ (.A(_122_),
    .B(_123_),
    .Y(_124_));
 sky130_fd_sc_hd__a21boi_1 _157_ (.A1(net17),
    .A2(_123_),
    .B1_N(_122_),
    .Y(_125_));
 sky130_fd_sc_hd__nand2_1 _158_ (.A(net7),
    .B(net30),
    .Y(_126_));
 sky130_fd_sc_hd__or2_1 _159_ (.A(net7),
    .B(net30),
    .X(_127_));
 sky130_fd_sc_hd__nand2_1 _160_ (.A(_126_),
    .B(_127_),
    .Y(_128_));
 sky130_fd_sc_hd__a21boi_1 _161_ (.A1(net16),
    .A2(_127_),
    .B1_N(_126_),
    .Y(_129_));
 sky130_fd_sc_hd__xor2_1 _162_ (.A(net17),
    .B(_124_),
    .X(_130_));
 sky130_fd_sc_hd__or2_1 _163_ (.A(_129_),
    .B(_130_),
    .X(_131_));
 sky130_fd_sc_hd__xor2_1 _164_ (.A(_129_),
    .B(_130_),
    .X(_132_));
 sky130_fd_sc_hd__nand2_1 _165_ (.A(net26),
    .B(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__nand2_1 _166_ (.A(_131_),
    .B(_133_),
    .Y(_134_));
 sky130_fd_sc_hd__a21o_1 _167_ (.A1(_131_),
    .A2(_133_),
    .B1(_125_),
    .X(_135_));
 sky130_fd_sc_hd__xor2_1 _168_ (.A(_125_),
    .B(_134_),
    .X(_136_));
 sky130_fd_sc_hd__or2_1 _169_ (.A(net26),
    .B(_132_),
    .X(_137_));
 sky130_fd_sc_hd__nand2_1 _170_ (.A(_133_),
    .B(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__xor2_1 _171_ (.A(net16),
    .B(_128_),
    .X(_139_));
 sky130_fd_sc_hd__nand2_1 _172_ (.A(net6),
    .B(net29),
    .Y(_140_));
 sky130_fd_sc_hd__or2_1 _173_ (.A(net6),
    .B(net29),
    .X(_141_));
 sky130_fd_sc_hd__nand2_1 _174_ (.A(_140_),
    .B(_141_),
    .Y(_142_));
 sky130_fd_sc_hd__a21boi_1 _175_ (.A1(net15),
    .A2(_141_),
    .B1_N(_140_),
    .Y(_143_));
 sky130_fd_sc_hd__or2_1 _176_ (.A(_139_),
    .B(_143_),
    .X(_144_));
 sky130_fd_sc_hd__xnor2_1 _177_ (.A(_139_),
    .B(_143_),
    .Y(_022_));
 sky130_fd_sc_hd__or2_1 _178_ (.A(_119_),
    .B(_022_),
    .X(_023_));
 sky130_fd_sc_hd__nand3_1 _179_ (.A(_138_),
    .B(_144_),
    .C(_023_),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _180_ (.A(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__xnor2_1 _181_ (.A(_119_),
    .B(_022_),
    .Y(_026_));
 sky130_fd_sc_hd__xor2_1 _182_ (.A(net15),
    .B(_142_),
    .X(_027_));
 sky130_fd_sc_hd__and2_1 _183_ (.A(net5),
    .B(net28),
    .X(_028_));
 sky130_fd_sc_hd__xor2_1 _184_ (.A(net5),
    .B(net28),
    .X(_029_));
 sky130_fd_sc_hd__a21oi_1 _185_ (.A1(net14),
    .A2(_029_),
    .B1(_028_),
    .Y(_030_));
 sky130_fd_sc_hd__nor2_1 _186_ (.A(_027_),
    .B(_030_),
    .Y(_031_));
 sky130_fd_sc_hd__xnor2_1 _187_ (.A(_027_),
    .B(_030_),
    .Y(_032_));
 sky130_fd_sc_hd__nor2_1 _188_ (.A(_118_),
    .B(_032_),
    .Y(_033_));
 sky130_fd_sc_hd__nor2_1 _189_ (.A(_031_),
    .B(_033_),
    .Y(_034_));
 sky130_fd_sc_hd__o21ba_1 _190_ (.A1(_031_),
    .A2(_033_),
    .B1_N(_026_),
    .X(_035_));
 sky130_fd_sc_hd__inv_2 _191_ (.A(_035_),
    .Y(_036_));
 sky130_fd_sc_hd__xnor2_1 _192_ (.A(_026_),
    .B(_034_),
    .Y(_037_));
 sky130_fd_sc_hd__xnor2_1 _193_ (.A(_118_),
    .B(_032_),
    .Y(_038_));
 sky130_fd_sc_hd__xnor2_1 _194_ (.A(net14),
    .B(_029_),
    .Y(_039_));
 sky130_fd_sc_hd__and2_1 _195_ (.A(net4),
    .B(net27),
    .X(_040_));
 sky130_fd_sc_hd__xor2_1 _196_ (.A(net4),
    .B(net27),
    .X(_041_));
 sky130_fd_sc_hd__a21oi_1 _197_ (.A1(net12),
    .A2(_041_),
    .B1(_040_),
    .Y(_042_));
 sky130_fd_sc_hd__or2_1 _198_ (.A(_039_),
    .B(_042_),
    .X(_043_));
 sky130_fd_sc_hd__xnor2_1 _199_ (.A(_039_),
    .B(_042_),
    .Y(_044_));
 sky130_fd_sc_hd__or2_1 _200_ (.A(_117_),
    .B(_044_),
    .X(_045_));
 sky130_fd_sc_hd__and3_1 _201_ (.A(_038_),
    .B(_043_),
    .C(_045_),
    .X(_046_));
 sky130_fd_sc_hd__xnor2_1 _202_ (.A(_117_),
    .B(_044_),
    .Y(_047_));
 sky130_fd_sc_hd__xnor2_1 _203_ (.A(net12),
    .B(_041_),
    .Y(_048_));
 sky130_fd_sc_hd__and2_1 _204_ (.A(net3),
    .B(net24),
    .X(_049_));
 sky130_fd_sc_hd__xor2_1 _205_ (.A(net3),
    .B(net24),
    .X(_050_));
 sky130_fd_sc_hd__a21oi_1 _206_ (.A1(net11),
    .A2(_050_),
    .B1(_049_),
    .Y(_051_));
 sky130_fd_sc_hd__nor2_1 _207_ (.A(_048_),
    .B(_051_),
    .Y(_052_));
 sky130_fd_sc_hd__xnor2_1 _208_ (.A(_048_),
    .B(_051_),
    .Y(_053_));
 sky130_fd_sc_hd__nor2_1 _209_ (.A(_116_),
    .B(_053_),
    .Y(_054_));
 sky130_fd_sc_hd__nor2_1 _210_ (.A(_052_),
    .B(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__o21ba_1 _211_ (.A1(_052_),
    .A2(_054_),
    .B1_N(_047_),
    .X(_056_));
 sky130_fd_sc_hd__inv_2 _212_ (.A(_056_),
    .Y(_057_));
 sky130_fd_sc_hd__xnor2_1 _213_ (.A(_047_),
    .B(_055_),
    .Y(_058_));
 sky130_fd_sc_hd__xnor2_1 _214_ (.A(net11),
    .B(_050_),
    .Y(_059_));
 sky130_fd_sc_hd__and2_1 _215_ (.A(net33),
    .B(net13),
    .X(_060_));
 sky130_fd_sc_hd__xor2_1 _216_ (.A(net33),
    .B(net13),
    .X(_061_));
 sky130_fd_sc_hd__a21oi_1 _217_ (.A1(net10),
    .A2(_061_),
    .B1(_060_),
    .Y(_062_));
 sky130_fd_sc_hd__or2_1 _218_ (.A(_059_),
    .B(_062_),
    .X(_063_));
 sky130_fd_sc_hd__xnor2_1 _219_ (.A(_059_),
    .B(_062_),
    .Y(_064_));
 sky130_fd_sc_hd__or2_1 _220_ (.A(_115_),
    .B(_064_),
    .X(_065_));
 sky130_fd_sc_hd__xnor2_1 _221_ (.A(_116_),
    .B(_053_),
    .Y(_066_));
 sky130_fd_sc_hd__and3_1 _222_ (.A(_063_),
    .B(_065_),
    .C(_066_),
    .X(_067_));
 sky130_fd_sc_hd__a21o_1 _223_ (.A1(_063_),
    .A2(_065_),
    .B1(_066_),
    .X(_068_));
 sky130_fd_sc_hd__xnor2_1 _224_ (.A(_115_),
    .B(_064_),
    .Y(_069_));
 sky130_fd_sc_hd__nand2_1 _225_ (.A(net32),
    .B(net2),
    .Y(_070_));
 sky130_fd_sc_hd__or2_1 _226_ (.A(net32),
    .B(net2),
    .X(_071_));
 sky130_fd_sc_hd__nand2_1 _227_ (.A(_070_),
    .B(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__a21boi_1 _228_ (.A1(net9),
    .A2(_071_),
    .B1_N(_070_),
    .Y(_073_));
 sky130_fd_sc_hd__xnor2_1 _229_ (.A(net10),
    .B(_061_),
    .Y(_074_));
 sky130_fd_sc_hd__nor2_1 _230_ (.A(_073_),
    .B(_074_),
    .Y(_075_));
 sky130_fd_sc_hd__xor2_1 _231_ (.A(_073_),
    .B(_074_),
    .X(_076_));
 sky130_fd_sc_hd__a21o_1 _232_ (.A1(net19),
    .A2(_076_),
    .B1(_075_),
    .X(_077_));
 sky130_fd_sc_hd__nand2b_1 _233_ (.A_N(_069_),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__xor2_1 _234_ (.A(_069_),
    .B(_077_),
    .X(_079_));
 sky130_fd_sc_hd__xor2_1 _235_ (.A(net9),
    .B(_072_),
    .X(_080_));
 sky130_fd_sc_hd__or2_1 _236_ (.A(_114_),
    .B(_080_),
    .X(_081_));
 sky130_fd_sc_hd__xnor2_1 _237_ (.A(net19),
    .B(_076_),
    .Y(_082_));
 sky130_fd_sc_hd__or2_1 _238_ (.A(_081_),
    .B(_082_),
    .X(_083_));
 sky130_fd_sc_hd__or2_1 _239_ (.A(_079_),
    .B(_083_),
    .X(_084_));
 sky130_fd_sc_hd__nand2_1 _240_ (.A(_078_),
    .B(_084_),
    .Y(_085_));
 sky130_fd_sc_hd__o211a_1 _241_ (.A1(_079_),
    .A2(_083_),
    .B1(_068_),
    .C1(_078_),
    .X(_086_));
 sky130_fd_sc_hd__nand2b_1 _242_ (.A_N(_067_),
    .B(_068_),
    .Y(_087_));
 sky130_fd_sc_hd__or3_1 _243_ (.A(_058_),
    .B(_067_),
    .C(_086_),
    .X(_088_));
 sky130_fd_sc_hd__a21o_1 _244_ (.A1(_043_),
    .A2(_045_),
    .B1(_038_),
    .X(_089_));
 sky130_fd_sc_hd__o311a_1 _245_ (.A1(_058_),
    .A2(_067_),
    .A3(_086_),
    .B1(_089_),
    .C1(_057_),
    .X(_090_));
 sky130_fd_sc_hd__nand2b_1 _246_ (.A_N(_046_),
    .B(_089_),
    .Y(_091_));
 sky130_fd_sc_hd__or3_1 _247_ (.A(_037_),
    .B(_046_),
    .C(_090_),
    .X(_092_));
 sky130_fd_sc_hd__a21o_1 _248_ (.A1(_144_),
    .A2(_023_),
    .B1(_138_),
    .X(_093_));
 sky130_fd_sc_hd__o311a_1 _249_ (.A1(_037_),
    .A2(_046_),
    .A3(_090_),
    .B1(_093_),
    .C1(_036_),
    .X(_094_));
 sky130_fd_sc_hd__nand2_1 _250_ (.A(_024_),
    .B(_093_),
    .Y(_095_));
 sky130_fd_sc_hd__or3_1 _251_ (.A(_136_),
    .B(_025_),
    .C(_094_),
    .X(_096_));
 sky130_fd_sc_hd__a31oi_1 _252_ (.A1(net47),
    .A2(_135_),
    .A3(_096_),
    .B1(_121_),
    .Y(_021_));
 sky130_fd_sc_hd__o21ai_1 _253_ (.A1(_025_),
    .A2(_094_),
    .B1(_136_),
    .Y(_097_));
 sky130_fd_sc_hd__and2b_1 _254_ (.A_N(net47),
    .B(net77),
    .X(_098_));
 sky130_fd_sc_hd__a31o_1 _255_ (.A1(net47),
    .A2(_096_),
    .A3(_097_),
    .B1(_098_),
    .X(_020_));
 sky130_fd_sc_hd__o31a_1 _256_ (.A1(_037_),
    .A2(_046_),
    .A3(_090_),
    .B1(_036_),
    .X(_099_));
 sky130_fd_sc_hd__xor2_1 _257_ (.A(_095_),
    .B(_099_),
    .X(_100_));
 sky130_fd_sc_hd__mux2_1 _258_ (.A0(net75),
    .A1(_100_),
    .S(net47),
    .X(_019_));
 sky130_fd_sc_hd__and2b_1 _259_ (.A_N(net47),
    .B(net41),
    .X(_101_));
 sky130_fd_sc_hd__o21ai_1 _260_ (.A1(_046_),
    .A2(_090_),
    .B1(_037_),
    .Y(_102_));
 sky130_fd_sc_hd__a31o_1 _261_ (.A1(net47),
    .A2(_092_),
    .A3(_102_),
    .B1(_101_),
    .X(_018_));
 sky130_fd_sc_hd__nand2_1 _262_ (.A(_057_),
    .B(_088_),
    .Y(_103_));
 sky130_fd_sc_hd__xnor2_1 _263_ (.A(_091_),
    .B(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__mux2_1 _264_ (.A0(net72),
    .A1(_104_),
    .S(net46),
    .X(_017_));
 sky130_fd_sc_hd__and2b_1 _265_ (.A_N(net46),
    .B(net39),
    .X(_105_));
 sky130_fd_sc_hd__o21ai_1 _266_ (.A1(_067_),
    .A2(_086_),
    .B1(_058_),
    .Y(_106_));
 sky130_fd_sc_hd__a31o_1 _267_ (.A1(net46),
    .A2(_088_),
    .A3(_106_),
    .B1(_105_),
    .X(_016_));
 sky130_fd_sc_hd__xnor2_1 _268_ (.A(_085_),
    .B(_087_),
    .Y(_107_));
 sky130_fd_sc_hd__mux2_1 _269_ (.A0(net74),
    .A1(_107_),
    .S(net46),
    .X(_015_));
 sky130_fd_sc_hd__and2b_1 _270_ (.A_N(net46),
    .B(net37),
    .X(_108_));
 sky130_fd_sc_hd__nand2_1 _271_ (.A(_079_),
    .B(_083_),
    .Y(_109_));
 sky130_fd_sc_hd__a31o_1 _272_ (.A1(net46),
    .A2(_084_),
    .A3(_109_),
    .B1(_108_),
    .X(_014_));
 sky130_fd_sc_hd__nand2_1 _273_ (.A(_081_),
    .B(_082_),
    .Y(_110_));
 sky130_fd_sc_hd__and2b_1 _274_ (.A_N(net46),
    .B(net36),
    .X(_111_));
 sky130_fd_sc_hd__a31o_1 _275_ (.A1(net46),
    .A2(_083_),
    .A3(_110_),
    .B1(_111_),
    .X(_013_));
 sky130_fd_sc_hd__and2b_1 _276_ (.A_N(net46),
    .B(net76),
    .X(_112_));
 sky130_fd_sc_hd__nand2_1 _277_ (.A(_114_),
    .B(_080_),
    .Y(_113_));
 sky130_fd_sc_hd__a31o_1 _278_ (.A1(net46),
    .A2(_081_),
    .A3(_113_),
    .B1(_112_),
    .X(_012_));
 sky130_fd_sc_hd__inv_2 _279_ (.A(net48),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _280_ (.A(net48),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _281_ (.A(net48),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _282_ (.A(net48),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _283_ (.A(net48),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _284_ (.A(net48),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _285_ (.A(net48),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _286_ (.A(net48),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _287_ (.A(net48),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _288_ (.A(net1),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _289_ (.A(net1),
    .Y(_011_));
 sky130_fd_sc_hd__dfrtp_1 _290_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(_012_),
    .RESET_B(_000_),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_1 _291_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(_013_),
    .RESET_B(_001_),
    .Q(net36));
 sky130_fd_sc_hd__dfrtp_1 _292_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(_014_),
    .RESET_B(_002_),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_1 _293_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(_015_),
    .RESET_B(_003_),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_1 _294_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(_016_),
    .RESET_B(_004_),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_1 _295_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(_017_),
    .RESET_B(_005_),
    .Q(net40));
 sky130_fd_sc_hd__dfrtp_1 _296_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(_018_),
    .RESET_B(_006_),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _297_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(_019_),
    .RESET_B(_007_),
    .Q(net42));
 sky130_fd_sc_hd__dfrtp_1 _298_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(_020_),
    .RESET_B(_008_),
    .Q(net43));
 sky130_fd_sc_hd__dfrtp_1 _299_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(_021_),
    .RESET_B(_009_),
    .Q(net44));
 sky130_fd_sc_hd__dfrtp_1 _300_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(net71),
    .RESET_B(_010_),
    .Q(net45));
 sky130_fd_sc_hd__dfrtp_1 _301_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(net34),
    .RESET_B(_011_),
    .Q(state));
 sky130_fd_sc_hd__conb_1 accelerator_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 accelerator_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 accelerator_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 accelerator_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 accelerator_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 accelerator_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 accelerator_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 accelerator_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 accelerator_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 accelerator_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 accelerator_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 accelerator_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 accelerator_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 accelerator_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 accelerator_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 accelerator_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 accelerator_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 accelerator_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 accelerator_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 accelerator_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 accelerator_70 (.LO(net70));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_87 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(arst_i),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(data_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(data_in[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(data_in[11]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(data_in[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(data_in[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(data_in[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(data_in[15]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(data_in[16]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(data_in[17]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(data_in[18]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(data_in[19]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(data_in[1]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(data_in[20]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(data_in[21]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(data_in[22]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(data_in[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(data_in[24]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(data_in[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(data_in[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(data_in[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(data_in[28]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(data_in[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(data_in[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(data_in[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(data_in[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(data_in[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(data_in[4]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(data_in[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(data_in[6]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(data_in[7]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(data_in[8]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(data_in[9]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(start),
    .X(net34));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(data_out[0]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(data_out[1]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(data_out[2]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(data_out[3]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(data_out[4]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(data_out[5]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(data_out[6]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(data_out[7]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(data_out[8]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(data_out[9]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(done));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(_120_),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(_120_),
    .X(net47));
 sky130_fd_sc_hd__buf_4 fanout48 (.A(net1),
    .X(net48));
 sky130_fd_sc_hd__conb_1 accelerator_49 (.LO(net49));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_1_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_1_1__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload0 (.A(clknet_1_0__leaf_clk_i));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(state),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net40),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net44),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net38),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net42),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net35),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net43),
    .X(net77));
 sky130_fd_sc_hd__decap_4 FILLER_0_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_113 ();
 assign data_out[10] = net49;
 assign data_out[11] = net50;
 assign data_out[12] = net51;
 assign data_out[13] = net52;
 assign data_out[14] = net53;
 assign data_out[15] = net54;
 assign data_out[16] = net55;
 assign data_out[17] = net56;
 assign data_out[18] = net57;
 assign data_out[19] = net58;
 assign data_out[20] = net59;
 assign data_out[21] = net60;
 assign data_out[22] = net61;
 assign data_out[23] = net62;
 assign data_out[24] = net63;
 assign data_out[25] = net64;
 assign data_out[26] = net65;
 assign data_out[27] = net66;
 assign data_out[28] = net67;
 assign data_out[29] = net68;
 assign data_out[30] = net69;
 assign data_out[31] = net70;
endmodule
