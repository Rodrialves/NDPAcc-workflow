`define ADDR_BUS_W 24
`define FE_ADDR_W 22
`define FE_DATA_W 32
`define BE_DATA_W 64
`define BE_ADDR_W 24
`define BE_STRB_W 8
`define FE_STRB_W 4
`define FIFO_DEPTH 16
